LIBRARY IEEE;
LIBRARY work;
USE work.MyPackage.all;

ENTITY TESTBENCH IS
END ENTITY;

ARCHITECTURE RTL OF TESTBENCH IS

	SIGNAL S_A      : INTEGER := 10;
	SIGNAL S_B      : INTEGER := 5;
	SIGNAL S_OP     : BIT_VECTOR (1 DOWNTO 0);
	SIGNAL S_OUTPUT : INTEGER;
	
BEGIN

    ALU_0 : ALU
	 PORT MAP (
		IN_A => S_A,
		IN_B => S_B,
		OP => S_OP,
		OUTPUT => S_OUTPUT
	);

	S_OP <= "00" AFTER 0ns, "01" AFTER 40ns, "10" AFTER 80ns, "11" AFTER 120ns;
		  
END ARCHITECTURE;